library verilog;
use verilog.vl_types.all;
entity SignExtend26_vlg_vec_tst is
end SignExtend26_vlg_vec_tst;
