library verilog;
use verilog.vl_types.all;
entity prueba1_vlg_vec_tst is
end prueba1_vlg_vec_tst;
