library verilog;
use verilog.vl_types.all;
entity uControl_vlg_vec_tst is
end uControl_vlg_vec_tst;
