library verilog;
use verilog.vl_types.all;
entity pruebaControl_vlg_vec_tst is
end pruebaControl_vlg_vec_tst;
