library verilog;
use verilog.vl_types.all;
entity InstructionReg_vlg_vec_tst is
end InstructionReg_vlg_vec_tst;
