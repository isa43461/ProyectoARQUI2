library verilog;
use verilog.vl_types.all;
entity prueba3_vlg_vec_tst is
end prueba3_vlg_vec_tst;
