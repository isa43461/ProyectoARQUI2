library verilog;
use verilog.vl_types.all;
entity prueba2_vlg_vec_tst is
end prueba2_vlg_vec_tst;
