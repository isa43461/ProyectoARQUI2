library verilog;
use verilog.vl_types.all;
entity Alu_vlg_vec_tst is
end Alu_vlg_vec_tst;
