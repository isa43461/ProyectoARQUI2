library verilog;
use verilog.vl_types.all;
entity RegFile_vlg_vec_tst is
end RegFile_vlg_vec_tst;
