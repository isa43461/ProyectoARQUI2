library verilog;
use verilog.vl_types.all;
entity AluControl_vlg_vec_tst is
end AluControl_vlg_vec_tst;
